module and32(out, in1, in2);
    input [31:0] in1, in2;
    output [31:0] out;
    and n0(out[0], in1[0], in2[0]);
    and n1(out[1], in1[1], in2[1]);
    and n2(out[2], in1[2], in2[2]);
    and n3(out[3], in1[3], in2[3]);
    and n4(out[4], in1[4], in2[4]);
    and n5(out[5], in1[5], in2[5]);
    and n6(out[6], in1[6], in2[6]);
    and n7(out[7], in1[7], in2[7]);

    and n8(out[8], in1[8], in2[8]);
    and n9(out[9], in1[9], in2[9]);
    and n10(out[10], in1[10], in2[10]);
    and n11(out[11], in1[11], in2[11]);
    and n12(out[12], in1[12], in2[12]);
    and n13(out[13], in1[13], in2[13]);
    and n14(out[14], in1[14], in2[14]);
    and n15(out[15], in1[15], in2[15]);

    and n16(out[16], in1[16], in2[16]);
    and n17(out[17], in1[17], in2[17]);
    and n18(out[18], in1[18], in2[18]);
    and n19(out[19], in1[19], in2[19]);
    and n20(out[20], in1[20], in2[20]);
    and n21(out[21], in1[21], in2[21]);
    and n22(out[22], in1[22], in2[22]);
    and n23(out[23], in1[23], in2[23]);

    and n24(out[24], in1[24], in2[24]);
    and n25(out[25], in1[25], in2[25]);
    and n26(out[26], in1[26], in2[26]);
    and n27(out[27], in1[27], in2[27]);
    and n28(out[28], in1[28], in2[28]);
    and n29(out[29], in1[29], in2[29]);
    and n30(out[30], in1[30], in2[30]);
    and n31(out[31], in1[31], in2[31]);
endmodule